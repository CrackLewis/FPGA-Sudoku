`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/01/02 20:46:24
// Design Name: 
// Module Name: NumberLattice
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module NumberLattice(
        number, lattice
    );
    input [3:0] number;
    output [120:0] lattice;

    wire [9:0] nums;
    assign nums[0] = (number == 4'd0);
    assign nums[1] = (number == 4'd1);
    assign nums[2] = (number == 4'd2);
    assign nums[3] = (number == 4'd3);
    assign nums[4] = (number == 4'd4);
    assign nums[5] = (number == 4'd5);
    assign nums[6] = (number == 4'd6);
    assign nums[7] = (number == 4'd7);
    assign nums[8] = (number == 4'd8);
    assign nums[9] = (number == 4'd9);
    // the following lattice is auto-generated by external programs.
    assign lattice[0] = 0;
    assign lattice[1] = 0;
    assign lattice[2] = 0;
    assign lattice[3] = 0;
    assign lattice[4] = 0;
    assign lattice[5] = 0;
    assign lattice[6] = 0;
    assign lattice[7] = 0;
    assign lattice[8] = 0;
    assign lattice[9] = 0;
    assign lattice[10] = 0;
    assign lattice[11] = 0;
    assign lattice[12] = 0;
    assign lattice[13] = nums[5] | nums[7];
    assign lattice[14] = nums[2] | nums[3] | nums[5] | nums[6] | nums[7] | nums[8] | nums[9];
    assign lattice[15] = nums[2] | nums[3] | nums[5] | nums[6] | nums[7] | nums[8] | nums[9];
    assign lattice[16] = nums[1] | nums[2] | nums[3] | nums[4] | nums[5] | nums[6] | nums[7] | nums[8] | nums[9];
    assign lattice[17] = nums[1] | nums[2] | nums[3] | nums[4] | nums[5] | nums[6] | nums[7] | nums[8] | nums[9];
    assign lattice[18] = nums[2] | nums[3] | nums[5] | nums[6] | nums[7] | nums[8] | nums[9];
    assign lattice[19] = nums[5] | nums[7];
    assign lattice[20] = 0;
    assign lattice[21] = 0;
    assign lattice[22] = 0;
    assign lattice[23] = 0;
    assign lattice[24] = nums[2] | nums[3] | nums[5] | nums[6] | nums[8] | nums[9];
    assign lattice[25] = 0;
    assign lattice[26] = nums[1] | nums[4];
    assign lattice[27] = 0;
    assign lattice[28] = nums[1] | nums[4];
    assign lattice[29] = 0;
    assign lattice[30] = nums[2] | nums[3] | nums[6] | nums[7] | nums[8] | nums[9];
    assign lattice[31] = 0;
    assign lattice[32] = 0;
    assign lattice[33] = 0;
    assign lattice[34] = 0;
    assign lattice[35] = nums[5] | nums[6] | nums[8] | nums[9];
    assign lattice[36] = nums[1];
    assign lattice[37] = nums[4];
    assign lattice[38] = 0;
    assign lattice[39] = nums[1] | nums[4];
    assign lattice[40] = nums[7];
    assign lattice[41] = nums[2] | nums[3] | nums[8] | nums[9];
    assign lattice[42] = 0;
    assign lattice[43] = 0;
    assign lattice[44] = 0;
    assign lattice[45] = 0;
    assign lattice[46] = nums[5] | nums[6] | nums[9];
    assign lattice[47] = nums[4] | nums[5] | nums[8];
    assign lattice[48] = nums[5] | nums[8];
    assign lattice[49] = nums[5] | nums[8];
    assign lattice[50] = nums[1] | nums[4] | nums[5] | nums[8];
    assign lattice[51] = nums[5] | nums[7] | nums[8];
    assign lattice[52] = nums[2] | nums[3] | nums[9];
    assign lattice[53] = 0;
    assign lattice[54] = 0;
    assign lattice[55] = 0;
    assign lattice[56] = 0;
    assign lattice[57] = nums[4] | nums[6] | nums[8];
    assign lattice[58] = nums[6] | nums[9];
    assign lattice[59] = nums[3] | nums[6] | nums[9];
    assign lattice[60] = nums[3] | nums[6] | nums[9];
    assign lattice[61] = nums[1] | nums[2] | nums[3] | nums[4] | nums[6] | nums[7] | nums[9];
    assign lattice[62] = nums[2] | nums[3] | nums[6] | nums[9];
    assign lattice[63] = nums[5] | nums[8] | nums[9];
    assign lattice[64] = 0;
    assign lattice[65] = 0;
    assign lattice[66] = 0;
    assign lattice[67] = 0;
    assign lattice[68] = nums[4] | nums[6] | nums[8];
    assign lattice[69] = nums[4];
    assign lattice[70] = nums[2] | nums[4];
    assign lattice[71] = nums[2] | nums[4];
    assign lattice[72] = nums[1] | nums[4] | nums[7];
    assign lattice[73] = nums[4];
    assign lattice[74] = nums[3] | nums[4] | nums[5] | nums[6] | nums[8] | nums[9];
    assign lattice[75] = 0;
    assign lattice[76] = 0;
    assign lattice[77] = 0;
    assign lattice[78] = 0;
    assign lattice[79] = nums[6] | nums[8];
    assign lattice[80] = nums[2];
    assign lattice[81] = 0;
    assign lattice[82] = nums[7];
    assign lattice[83] = nums[1] | nums[4];
    assign lattice[84] = 0;
    assign lattice[85] = nums[3] | nums[5] | nums[6] | nums[8] | nums[9];
    assign lattice[86] = 0;
    assign lattice[87] = 0;
    assign lattice[88] = 0;
    assign lattice[89] = 0;
    assign lattice[90] = nums[2] | nums[3] | nums[5] | nums[6] | nums[8];
    assign lattice[91] = 0;
    assign lattice[92] = 0;
    assign lattice[93] = nums[7];
    assign lattice[94] = nums[1] | nums[4];
    assign lattice[95] = nums[9];
    assign lattice[96] = nums[3] | nums[5] | nums[6] | nums[8];
    assign lattice[97] = 0;
    assign lattice[98] = 0;
    assign lattice[99] = 0;
    assign lattice[100] = 0;
    assign lattice[101] = nums[1] | nums[2];
    assign lattice[102] = nums[1] | nums[2] | nums[3] | nums[5] | nums[6] | nums[8];
    assign lattice[103] = nums[1] | nums[2] | nums[3] | nums[5] | nums[6] | nums[8] | nums[9];
    assign lattice[104] = nums[1] | nums[2] | nums[3] | nums[5] | nums[6] | nums[7] | nums[8] | nums[9];
    assign lattice[105] = nums[1] | nums[2] | nums[3] | nums[4] | nums[5] | nums[6] | nums[8] | nums[9];
    assign lattice[106] = nums[1] | nums[2] | nums[3] | nums[5] | nums[6] | nums[8];
    assign lattice[107] = nums[1] | nums[2];
    assign lattice[108] = 0;
    assign lattice[109] = 0;
    assign lattice[110] = 0;
    assign lattice[111] = 0;
    assign lattice[112] = 0;
    assign lattice[113] = 0;
    assign lattice[114] = 0;
    assign lattice[115] = 0;
    assign lattice[116] = 0;
    assign lattice[117] = 0;
    assign lattice[118] = 0;
    assign lattice[119] = 0;
    assign lattice[120] = 0;
endmodule
