`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/01/01 15:22:41
// Design Name: 
// Module Name: GameTemplate
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module GameTemplate(
        sig_new, seed,
        template_map
    );
    input sig_new;
    input [31:0] seed;
    output [323:0] template_map;

    wire [323:0] base [127:0];
    assign base[0]  = 324'b001010011000000101000110001101010111000101100101001101110010010010001001001101110100010110001001000100100110010000100001011010010011010101111000011010000011010001010111100100010010100101010111001000011000011000110100100000110010100101100001011101000101011101000110100000110101001010010001010100011001011100100100100001100011;
    assign base[1]  = 324'b001110010101100001110010000101000110011000100001010101001001100000110111011101001000001100010110100100100101010101111001001001100100001100011000100001100100100100110001011101010010000100110010011110000101010001101001001001010111010010010011011010000001100100010011011001011000001001110100010010000110000100100111010110010011;
    assign base[2]  = 324'b011000100100001100010101100001111001000101110101001010011000010000110110001110001001010001110110001001010001010100011000011101000011011010010010011110010010010101100001001101001000010001100011100110000010011100010101100101000110100001010111000100100011001001010001011000110100100110000111100000110111000100101001010101100100;
    assign base[3]  = 324'b001100100001011110000100010110010110010001010110001100101001000110000111100101111000000101010110001101000010001010000111010110010011010001100001011000110100001000011000011101011001000110010101011001000111001000111000010100011001100000110010011001110100011101000010100101100101100000010011100001100011010001110001100100100101;
    assign base[4]  = 324'b100101100010001101000111010110000001000101000111100001100101001100101001100000110101000100101001011101100100010110000001001010010011011001000111001100100100011001111000000110010101011001111001010001010001001000111000001000010110010110000100100101110011011101011000100100110010010000010110010010010011011100010110100001010010;
    assign base[5]  = 324'b010110000011100101000010000101100111100100010111001110000110001001000101010001100010000101110101100100111000001010010110010100010111001110000100100001000101011000100011011100011001001101110001010010011000010100100110011000111000011101010001010010010010011100100100100000111001011001010001000101011001001001100100100001110011;
    assign base[6]  = 324'b001000011000011101100100001101011001010000110101001010011000000101110110100101110110010100010011010010000010011101010011011000100001100010010100100010010001010000110101001001100111011000100100100001111001010100010011001101100010000110000111100101000101010110000111100101000010011000110001000101001001001101010110011100101000;
    assign base[7]  = 324'b010000100101000100110111100101101000001100011000010001101001011100100101011110010110010100101000000100110100100000110100100100010010011001010111100101110001001101010110010010000010010101100010011110000100001110010001011001010011100001000001001001111001000110001001001001110011010101000110001001000111011010010101100000010011;
    assign base[8]  = 324'b001010001001011100110001010101000110001101010100011010001001011100100001011100010110001001010100100000111001010010010010100000010101001101100111010101100011010000100111100100011000000101111000100101100011010001010010100100100001001101001000011001110101011001000111010110010010000110000011100000110101000101110110001010010100;
    assign base[9]  = 324'b001001011001011001110011010000011000001100011000100100100100011001010111011001110100000101011000100100100011010000110010011110000001010110010110011101100001001010010101100000110100100010010101001101000110000101110010100101000011100000010010011101100101000110000110010100110111001001001001010100100111010001101001001110000001;
    assign base[10] = 324'b100100010111011000100101010000111000011010000101010000110111000100101001010000100011100100011000010101100111000101011000001101000110100101110010011101000010100001011001001100010110001110010110000101110010100001000101010101110100001010010011011010000001001001100001010110000100011110010011100000111001011101100001001001010100;
    assign base[11] = 324'b100100010100011000110111001001011000011000110101100110000010010000010111001001111000010001010001100100110110000101000011100001110110010100101001100000101001001100010101011001110100011101010110001010010100000110000011010010000010000101100011011110010101010110010001011101001000001101100010001101100111010100101001100001000001;
    assign base[12] = 324'b011110010100001001011000001100010110000110000011011001111001010100100100010101100010000100110100011110001001011001000111100000100001100100110101100100100101001101000111000101101000100000110001010110010110001001000111001000010110100110000101010001110011001101111001010001100010100001010001010001011000011100010011011010010010;
    assign base[13] = 324'b100110000001010001100011010100100111001101110100001000010101011010001001001001100101011110011000001100010100010000100110000101011001011100111000011101010011100001000110001010010001100000011001001101110010010001010110010110011000011000100111000101000011000100110111010110000100100101100010011001000010100100110001100001110101;
    assign base[14] = 324'b011100011001001101000101001010000110100000100011011101101001010100010100010101100100001010000001001101111001001101001000000100100111011010010101001010010111011001010100000100111000011001010001100010010011010000100111100100110101010001110010100001100001010010000010100100010110011101010011000101110110010100111000100101000010;
    assign base[15] = 324'b001010000011010100010100011010010111011001110100100100110010010100011000100100010101011101101000010000110010011110010010001101000101100001100001010000111000011010010001011100100101000101010110001010000111001101001001010100100001010001110110100110000011100001001001000101010011001001110110001101100111100000101001000101010100;
    assign base[16] = 324'b000100100111100001000110001110010101010100111000100100010111010001100010010010010110001000110101100000010111001001100011011110000100000101011001011100010100010101101001001000111000100001011001001100100001011101000110011010000101010001110011100100100001100101000010000101011000011001110011001101110001011010010010010110000100;
    assign base[17] = 324'b010110010100001101100001100001110010011100111000010000100101000101101001001000010110100010010111001101000101001100101001000101000110010110000111000110000111010100110010011010010100010001100101011110001001001000010011100101010010011000010100011100111000011001000011001001111000100101010001100001110001100101010011010000100110;
    assign base[18] = 324'b011110010110010100110100001010000001000100100011011010001001011101000101010001011000011100100001011010010011100000010101001110010110010001110010001101111001010000010010010101101000011001000010100001010111001100011001001010000100100101110011000101010110010100110111000101101000100100100100100101100001001001000101100000110111;
    assign base[19] = 324'b011100100001100101000110010110000011010110000100000100110111100100100110001110010110001001011000000101000111001000111000011000010101011110010100100100010111010000100011011001011000011001000101100001111001001000110001100001110011010101100010010000011001000101100010001110010100100001110101010001011001011110000001001101100010;
    assign base[20] = 324'b001010000110000101010100001101111001010000010011001001111001010110000110100101010111001110000110000101000010100000110100100100100001011001010111011000100001011101000101100010010011011110010101100001100011010000100001010101001001011000010111001000111000000101110010010000111000100101100101001101101000010110010010011100010100;
    assign base[21] = 324'b010001100101011100011000001110010010100010010111001100100101000101100100001100100001010001101001011101011000011100011000011001000011100100100101010101001001000110000010011000110111001000110110010110010111010010000001011010000010100101110100010100010011000101010100100000110110001001111001100101110011001001010001100001000110;
    assign base[22] = 324'b001001010100011001111000001100011001100100110110010100100001100001110100000101111000100100110100001001010110001110010001100001010110010000100111010001100111001100010010010110011000100000100101011101001001011000110001011000010010010010010011011110000101010110001001001001100111000101000011011101000011000110000101100101100010;
    assign base[23] = 324'b001000110100100101010001011010000111100110000101011100110110000100100100011001110001010000101000100100110101010101000011100010010111001000010110011100011001001001100101100001000011100001100010001100010100011101011001010000100110000101110011010110011000001110010111010110000010010001100001000101011000011001001001001101110010;
    assign base[24] = 324'b001110000010011101000001010101101001010100010110001010001001011101000011010010010111010101100011001010000001011001001000000110010010001101010111100101010001001101110110010000101000011100100011010001011000000110010110001000111001011000010100100001110101100001110100100100110101011000010010000101100101100000100111100100110100;
    assign base[25] = 324'b011000100101011100111000000110010100011101000001011001011001001100101000100010010011010000010010010101110110001000011001010101000011011010000111001110000110001010010111010001010001010101110100100001100001100100110010100101100010001110000100011100010101000101010111100100100110100001000011010000111000000101110101001001101001;
    assign base[26] = 324'b001001100100001110000001100101010111100100110101011100100100100000010110011100011000011010010101010000100011100001001001001001010110011100110001001101110110100000011001001001000101010100100001010000110111011010001001000101010010100101101000001101110100010010010011000101110010010101101000011010000111010101000011000110010010;
    assign base[27] = 324'b001100010100011000101000010101111001011100101000010010010101001101100001100101010110000101110011010000101000001001111001010100110001011010000100100001000001100101100111001000110101011000110101100001000010000110010111010110000010011100010110100101000011000110010011001010000100011101010110010001100111001101011001100000010010;
    assign base[28] = 324'b010100101000010000010011011110010110010010010001100001100111001001010011011100110110010110010010000110000100100101110101001100100110010000011000011010000010000101010100100100110111000101000011011110001001010101100010001000010100011000110101100001111001001101010111100101001000011000100001100001101001001001110001001101000101;
    assign base[29] = 324'b010101000011000110010010100001100111100001100001001101000111001001011001011100101001100001010110001101000001001001010100011100011000011010010011000110010110001000110101011110000100001110000111010001101001010100010010100100010010010110000011010001110110011000110101100101110100000100101000010001111000011000100001100100110101;
    assign base[30] = 324'b001001110110000110000101010010010011010100111000001010010100011000010111000110010100001101100111001010000101100100100001010001110011010101101000100001010011011000100001100101110100010001100111100001011001001100100001011001000010010100011000011100111001001100011001011101000010100001010110011110000101100100110110000101000010;
    assign base[31] = 324'b011001000111001010001001000101010011100001010010001101000001011010010111001110010001010101110110001001001000011110000101010010010010001100010110100100010100011101100011010110000010001001100011100000010101010001111001010101110110000100111000100100100100000100111000100100100100011101100101010000101001011001010111100000110001;
    assign base[32] = 324'b001000010100100001100101011110010011011010001001001001110011010101000001011101010011100101000001001001101000010100100111000100111001011010000100010010010001011001011000001101110010001101101000011100100100100100010101100001000110010110010010000100110111000101110010001110000110010001011001100100110101010000010111100000100110;
    assign base[33] = 324'b010000111001001010000101011101100001001000011000011100110110100101010100011101010110000110010100001010000011001110010001010000101000010101110110100001110101001101100001010010010010011001000010100101010111000100111000010100100011011000011001100001000111100101100100100001110010001100010101000110000111010101000011011000101001;
    assign base[34] = 324'b001000010101100100110100011110000110011110000011011000100001010101001001100101100100011110000101001000110001000100101001100001010110001101110100010101000110001001110011100100011000001101111000000101001001011000100101011010010010010000010111100001010011100000110001010110010010010001100111010001010111001101101000000110010010;
    assign base[35] = 324'b011001000101001010001001001100010111000101110011010001100101100000101001100110000010001100010111010101000110001001101001100001110011010001010001011101011000000101000110001010010011001100010100010110010010011001111000010000100111011000110001100110000101010110010110011100101000000100110100100000110001100101010100011101100010;
    assign base[36] = 324'b001001110110001101000101000110001001100000110001100100100110010101110100010101001001000101111000001100100110011000011000001000110111010010010101010010010101100001100001011100110010011100100011010110010100100001100001001101100111010000011001001001011000100101010100011110000010011000010011000110000010011001010011100101000111;
    assign base[37] = 324'b000101000011010110010010100001100111001010010111100001100011000101010100011001011000011100010100001000111001100001110001001000110101100101000110100100100101010010000110011100010011001101100100100101110001010110000010010110000110001100100111010010010001010000010010011001011001001101111000011100111001000101001000011000100101;
    assign base[38] = 324'b001001110100010100110001011010011000100000110001010001101001010100100111100101100101001001111000001100010100011101000010000110010011100001100101000110011000011001010111001001000011011001010011100000100100100101110001010100010111100110000010010000110110001100100110011101000101000110001001010010001001001100010110011101010010;
    assign base[39] = 324'b000100100111001110010101010001101000010101000011000110000110100101110010100101101000010000100111000100110101011000110001001001010100011110001001010010010101100001110001001100100110100001110010100101100011010101000001011100010110010101000010100010010011001110000100011000011001001001010111001001011001011100111000011000010100;
    assign base[40] = 324'b010000010110001000111001010101111000011100101000011001010100001100011001001110010101100000010111010000100110010101000001001110000010100101100111011001110011000110010101001010000100001010001001011101000110000100110101100001010111100100100001011001000011000100110100010101101000011110010010100101100010010001110011100001010001;
    assign base[41] = 324'b010000101000010110010001011001110011011110010101010001100011001010000001011000110001100000100111010010010101100001000110100100010010001101010111010101110010011000111000100100010100100100010011011101010100100000100110001110001001000101110110010101000010000101100100001010000101011100111001001001010111001101001001000101101000;
    assign base[42] = 324'b001110001001001000010100010101110110010000010111011001011000001100101001010100100110011110010011000101001000000110010101100000110111010001100010011001111000010000100101100100010011001001000011000101101001100001010111100001100010100101000001011100110101011101010100001110000110001010010001100100110001010101110010011010000100;
    assign base[43] = 324'b011010000010010000110111000110010101010001110101100100100001001110000110100100110001010110000110011101000010011100010011100001100100001001011001010101001001000101110010100001100011100000100110001101011001010000010111000101010111011001000011100100101000001101100100001010011000010101110001001010011000011100010101011000110100;
    assign base[44] = 324'b100001000010011001110001001110010101010100010011001001001001011010000111100101100111001110000101001001000001000101110101010001100010100000111001001110000100010110010111000101100010011000101001100000010011010101110100010010011000000100100110011101010011011100110001100101011000010000100110001001010110011100110100100100011000;
    assign base[45] = 324'b100001100001001000110100011101011001011100100101000101101001001110000100010010010011010101111000001001100001010110000111011000010011100101000010100100110100100000100111010100010110011000010010100101000101100000110111000101001001001101010010011001111000001001010110011110000001010010010011001101111000010010010110000100100101;
    assign base[46] = 324'b100000110010000110010101011001110100011101000001001001100011100010010101100101100101100001000111000100110010010000100011010100011000011101101001011000010111100100100100001101011000010110001001011100110110001001000001000101010110001110001001010000100111001010010100011001110001010110000011001101111000010001010010100100010110;
    assign base[47] = 324'b011010010100100000100001010100110111011100100011010001011001011010000001000110000101011001110011010000101001001001100001010110010111100001000011100101010111001110000100000101100010010000111000001000010110011110010101100001110110000100110010100101010100010100010010100101001000001101110110001101001001011101100101001000011000;
    assign base[48] = 324'b100100100110000100110100011110000101010001010001001001111000011010010011011110000011010110010110001000010100011001110100100100010101100000110010001110010010011010000111010001010001010100011000001101000010100101100111100000110111010001100001010100101001000101100101011100101001001101001000001001001001100001010011000101110110;
    assign base[49] = 324'b011001110011100000010010100101010100000110010010001101010100011110000110100001010100011101101001001100010010001101100001100101001000010100100111010101000111011000100001100010010011100100101000010101110011011001000001001000111001010010000111000101100101010010000110000100110101001001111001011100010101001010010110010000111000;
    assign base[50] = 324'b010100110001100001110100001001101001100101000010000100110110100001010111011101101000010100101001010000110001000101011001001001000111001110000110001001110110001100011000010110010100010010000011100101100101011100010010001100100101011110010001011001001000100000010100011001010010100101110011011010010111010010000011000100100101;
    assign base[51] = 324'b000100100110001101000101011110001001010101110011100010010110001001000001100110000100000101110010010100110110001110010101011010000111010000010010001001101000010001010001001110010111010000010111001000111001011001011000011100110001010100101000100101100100100001000010100101100011000101110101011001011001011100010100100000100011;
    assign base[52] = 324'b011100011000011000110100010110010010010100110010100010010111000101000110100101100100010100100001001110000111010001110011000101011001011000101000000110000110001101000010100101110101001010010101011110000110010000010011001100100001100101101000011101010100100001010111010000010011001001101001011001001001001001110101100000110001;
    assign base[53] = 324'b011110000001010101100100001100101001010100100100001110010001011010000111011010010011100001110010010100010100100101110010000110000011010001010110001101000110001001011001000101111000100000010101011001000111100100110010000101100111010000111000001010010101001001011000100100010110011101000011010000111001011100100101100001100001;
    assign base[54] = 324'b100101010110001110000100001000010111010000010111010110010010011000111000100000100011011101100001010010010101001001001001000101010110011110000011011000110101100001000111100100100001011110000001100100100011010101100100001101101000001001110101000101001001010110010100011000011000001101110010000101110010010000111001100001010110;
    assign base[55] = 324'b100000010101011100100100100101100011011110010011011010000001001001000101001001100100001101011001100001110001010001111001010100111000000100100110011000110001100101110010010110000100010100101000000101000110011100111001001101000111001010010101011000011000000101010010100001100011010010010111100110000110010000010111001101010010;
    assign base[56] = 324'b011101000010100101100011000110000101011000111001100000010101011100100100000110000101001001000111100100110110010100100110001110010001100001000111010001110011010110000110001000011001100010010001011100100100011001010011100101010100000101110010001101101000001001101000010000111001010101110001001100010111011001011000010010010010;
    assign base[57] = 324'b100001111001001001000011010100010110001101000101000101110110001010011000011000010010010110001001010001110011010100100011100101100001011110000100000110010111010000111000011000100101010010000110011100100101000100111001100101010100100000010010001101100111001001101000001101010111100101000001011100110001011010010100100001010010;
    assign base[58] = 324'b000100100110100001010111001101001001010001111001001100100001011010000101010110000011011001001001001000010111100100110100000101110110010100101000011000011000010110010010010001110011011101010010010010000011000110010110001101100111001000011000100101010100001010010101011100110100100001100001100001000001100101100101011100110010;
    assign base[59] = 324'b001001100001100100110100010110000111001101110101001001101000100100010100100010010100011101010001001001100011011001000010000101110101100000111001011101011001001110000010000101000110000100111000010010010110011100100101010100010011100001001001011001110010100110000111011000100011010001010001010000100110010100010111001110011000;
    assign base[60] = 324'b010110011000001101000001011100100110011100110110100100100101100001000001010000100001011001111000100101010011100001100111000101010100001000111001001001010011100010010110000101110100100100010100011100110010011010000101011001000101001000010111001110011000001110000010010001101001010100010111000101111001010110000011010001100010;
    assign base[61] = 324'b010000100001100101110101011000111000010101101001100000100011011100010100001101111000000101100100100100100101011100010011010010000110010110010010100101000010010100010111100001100011011010000101001000111001010001110001000110010100011101010010001110000110100001010110001110010001001001000111001000110111011001001000000101011001;
    assign base[62] = 324'b100000010110010101111001010000100011011101001001001100100001011010000101001001010011010010000110011110010001100110000001011101000011001001010110011000110101001010011000000101110100010000100111000101100101100000111001010101110010100100010100001101101000001101100100100001010010100100010111000110011000011000110111010101000010;
    assign base[63] = 324'b100000111001001001110110010101000001010001100111001101010001100000101001000101010010100010010100001101100111100110000101011000010111001000110100011000010011010000100101100101111000001001110100100110000011011000010101011101000110010100111001000110000010010100100001011101101000010010010011001110011000000101000010011101010110;
    assign base[64] = 324'b001010000011010001100111000101011001000101100111100110000101001001000011010001011001000100110010011110000110001101001000011100100110010110010001011100100001001101011001100001100100010110010110100001000001001101110010011000010100001001111000100100110101100000110010010110010100011000010111100101110101011000010011010000101000;
    assign base[65] = 324'b100101010100100000010111011000110010001100010110010001010010100010010111001001111000100100110110000101010100011001000001010100101001011110000011011110000010000101100011100101000101010100111001011101001000001000010110000110010101011001110100001100101000010000100111001110000001010101101001100001100011001010010101010001110001;
    assign base[66] = 324'b001001100001010101000111100100111000011101010100100100111000001001100001100000111001011000010010010001110101011001110101010010010011000110000010000110011000011100100110001101010100001101000010100001010001011110010110100110000110000101110100010100100011010100010011001010001001011001000111010000100111001101100101100000011001;
    assign base[67] = 324'b011000100001011110010100100000110101011110001001001101010110001001000001010000110101000100101000100101100111001010010100100000110101000101110110100001010110001000010111001110010100000101110011010001101001010100101000001100011000011001000010011101011001100101100010010101110001010010000011010101000111100110000011011000010010;
    assign base[68] = 324'b011100100110010001010011100100011000100001010100000110010010001101110110100100010011011101101000010101000010010010010101100001110001011000100011011001110001001000110101010010001001001000111000011001001001011101010001000101100111001110000100001010010101010101000010100100010110100000110111001110001001010100100111000101100100;
    assign base[69] = 324'b010000010111001100101000011010010101100001101001010101110001001000110100001100100101010010010110011100011000011100110001011001010010010010001001001010010110100001000011000101010111010101001000011100011001001100100110000101110010100110000100010101100011100101010011001001100111100001000001011010000100000100110101100101110010;
    assign base[70] = 324'b100100010100010101101000001100100111011000100111100101000011100000010101010110000011011100010010100101000110001101110110010001011001001010000001100001011001011000100001011100110100001001000001001110000111010101101001010000110101001010010110000101111000000101100010100001110101010010010011011110011000000100110100011001010010;
    assign base[71] = 324'b011000110010010101110100000110011000010001111001001010000001010101100011010100011000001101101001011101000010011100100011011000011000100101010100100101010110010000110010100000010111100001000001100101010111001100100110001110000100000110010110001001110101000101100101011100100011010010001001001010010111100001000101011000110001;
    assign base[72] = 324'b011000100111010010010011010100011000010100010100100001110010011000111001001110011000011001010001001001110100001001110001001101101000010010010101100001010011100100010100011101100010010001101001010100100111000110000011100110000101011101000110001100100001011100110010000110000101100101000110000101000110001000111001100001010111;
    assign base[73] = 324'b100101010111001100010100001010000110010010000001011001010010011100111001001001100011011110001001000101010100010100010100001000111000100101100111100000101001010101100111010000010011001101110110010010010001010100101000011110011000000100100011011001000101000100110101100101000110100001110010011001000010100001110101001110010001;
    assign base[74] = 324'b011100010100001101011000001010010110100000100101011010010100001100010111011010010011001001110001100001000101100100111000010001100111010100100001000101000010100110000101011001110011010101110110000100110010010010001001001001101001011101000011000101011000001110000001010100101001011101100100010001010111100000010110100100110010;
    assign base[75] = 324'b100000110110010110010111001000010100100101000111000101100010010110000011000100100101100000110100100101110110010001101000100100100011000101010111010100011001010001111000001101100010001101110010011001010001010010011000011010000001001001001001011100110101001001010011011100010110100001001001011110010100001110000101011000100001;
    assign base[76] = 324'b010000110110011100101001100000010101001000011000010000110101011001111001100101010111000101101000001101000010010110000010001101000111100101100001000101000011010110010110001010000111011001111001001010000001010100110100001110010100011000010010011101011000011100100001100001010011010010010110100001100101100101110100000100100011;
    assign base[77] = 324'b011101000101000100100011011010011000000100111000100101100100011100100101100101100010010101111000000100110100001110010111001010000001010001010110011000100100011100110101100000011001010110000001011001001001001001110011010001011001100000010010001101100111100000010110001101010111100101000010001001110011010010010110010110000001;
    assign base[78] = 324'b001000010100001101011000011010010111001101111001001001100001010101001000011010000101010010010111000100100011100101010010011001110011100000010100000101100111100001001001001000110101010000111000010100010010100101110110100001000001011100100110001101011001011100100110100100110101010010000001010110010011000110000100011101100010;
    assign base[79] = 324'b001100100100100101110110100001010001100010010110001101010001011100100100010100010111010000101000100100110110001001011001000101000111011010000011011001111000010110010011010000010010010000110001100001100010010101111001011101000101001000011001001101101000100110000010011000110101000101000111000101100011011110000100001010010101;
    assign base[80] = 324'b000110000110001001000111001110010101001101111001100001010001010000100110001001010100001101101001011100011000100001000001011010010010010100110111010101100010010001110011000110001001011110010011010100011000001001100100010000110101000110000110100101110010011000100111100100110101100001000001100100011000011100100100011001010011;
    assign base[81] = 324'b001010010101100000010110001101110100001101001000011101011001001001100001011101100001001001000011010110001001010100010100011000110010011110011000100100100011010001111000011000010101100001110110000110010101010000100011000100111001010101100111100001000010010010000111001100100001100101010110011001010010100110000100000100110111;
    assign base[82] = 324'b011110010001010010000101001001100011010001100011000100100111100001011001100001010010001101101001011101000001100100100101100001110011011000010100011010000111010101000001100100110010001100010100011010010010010110000111010101110110001000110100000110011000001000111000100100010110010001110101000101001001011101011000001100100110;
    assign base[83] = 324'b010101100001010001110010100000111001100110000010001101100101010000010111001101110100000110011000010100100110100000110101011001000111001010010001010010010110001010000001001101110101000100100111100101010011011001001000011101001001010100110110000110000010011000011000011100100100100101010011001001010011100000011001011101100100;
    assign base[84] = 324'b010101101000000101110010001110010100001000011001001101000101100001100111011100110100100010010110010100100001100101000111010101101000000100110010001110000010010000010111100101010110000101010110100100100011010001111000010000100001011101011001011010000011011010010011001010000100011100010101100001110101011000110001001001001001;
    assign base[85] = 324'b100110000100000101010011001001100111001000010101100101100111001101001000011101100011010000101000010110010001000110010110001010000101010001110011010001110010001100011001011010000101010100111000011101000110000100101001001100101001010101110100100000010110100001000111011000110001100101010010011001010001100010010010011100110100;
    assign base[86] = 324'b100000011001010101100011001001000111010001110011100000100001010101101001011000100101010001111001001100011000010110000001011000110100100101110010011101100010100110000101010000110001100100110100001000010111100001010110001110010110000101001000011100100101001001001000011101010110000110010011000101010111001110010010011010000100;
    assign base[87] = 324'b001001101000010100110111100100010100000101110100001010010110010110000011100101010011100000010100001001100111011000100111100110000001010000110101100000011001010001010011011100100110010000110101011101100010100010010001010110010001001101001000011001110010011101000110000100101001001101011000001110000010011001110101000101001001;
    assign base[88] = 324'b010000100110000110000011011110010101000101010011001010010111100001100100100101111000010001100101001000010011010100110111011001000010100110000001011010000001010100111001010001110010001010010100100001110001001101010110001101100010011101011000000101001001100000010101100100100100011000110111011101001001001100010110010100101000;
    assign base[89] = 324'b001101100100100101110101000100101000000110011000001000110110010101000111010101110010010010000001011000111001011000010111001100101000100101010100010010001001010101100111001000010011001001010011000101001001011110000110011101000110100001010010001110010001100100110101011000010100100001110010100000100001011110010011010001100101;
    assign base[90] = 324'b011100111001100000010010010101000110011000010100010110010111001100101000100001010010010000110110000110010111001110011000011101100100001001010001010000100111000101010011011010001001000101100101001010001001010001110011100110000001001101000101011101100010001001000011011001111000100100010101010101110110100100100001100000110100;
    assign base[91] = 324'b010100100001100110000111001101000110011100110110001001000001010110001001100001001001010100110110011100010010001010010111000101101000010001010011001100010101011110010100011000101000010001101000001101010010100101110001000101010010011001110011100010010100100110000011010000100101000101100111011001110100100000011001001000110101;
    assign base[92] = 324'b001101011001010000101000000101110110100001110001010100110110010010010010001001000110011110010001010110000011011101100101001010001001001101000001100100010010011001000011100001010111010010000011000101010111001001101001010100110100100101100010011100011000000110011000001101110100011000100101011000100111100000010101100100110100;
    assign base[93] = 324'b100100110001010010000110001001110101010110000010001100010111011001001001010001100111100100100101001100011000100000010100001001100011010110010111011100100011010110010001010010000110011010010101100001110100000100110010000101011001011101000010100001100011001001001000011000111001011101010001001101110110000101011000100100100100;
    assign base[94] = 324'b011010010001100001000010001101110101011101000101000100110110100100101000001110000010100101110101000101100100010101111000001100010100001010010110000101100011001001011001010010000111100100100100011010000111010100010011001001010111010010011000011000110001010000110110011100100001100001011001100000011001010101100011011101000010;
    assign base[95] = 324'b100001100011010000101001000101010111010001010111000100111000011000101001000100101001010101110110001101001000010100011000001110010010010001110110011001110010100001000101100100110001001110010100011000010111010110000010100100110110001010000100011100010101001001000101011101100001100010010011011110000001100101010011001001100100;
    assign base[96] = 324'b100001110101010000100110100100010011000110010010010100111000011101100100011001000011011100011001010100101000100101010001001110000010011001000111010000100111011001010001001110001001001110000110100101110100001001010001011100011001001001000101100000110110010100111000000101100111010010010010001001100100100010010011000101110101;
    assign base[97] = 324'b000100100110010001110011010110001001100001001001010100010010011000110111011100110101011010011000000101000010010110010111000110000110001100100100001001100001001101001001011101011000010010000011011100100101100100010110001101111000001001100001010010010101011000010010100101010100100001110011100101010100100000110111001001100001;
    assign base[98] = 324'b100100100011100001100101010001110001100001000101000100100111001101101001011000010111001101001001100000100101011101100100100100111000010100010010001110010001001001010110011110000100010110000010010001110001011010010011000101010110011110010100001000111000010000111001011010000010000101010111001001111000010100010011100101000110;
    assign base[99] = 324'b001100011000011101000101001001101001011100100100100101101000000100110101010110010110000100100011100001110100011000110010010010001001010100010111000101001001001001010111011010000011100001010111011000110001100101000010100101100101100001110100001100100001001001110011010100010110010010011000010010000001001110010010011101010110;
    assign base[100] = 324'b010100100001001110010110100001000111100001000011011100100001010101101001011010010111010110000100000100100011000101100100001001110101001110011000100101010010010000111000011001110001001101111000000101101001001001010100001000111001100001010111010000010110010010000110100100010010011100110101011100010101011001000011100110000010;
    assign base[101] = 324'b001001010100000101110011100101101000100000110110010010010101000101110010011110010001100001100010010000110101000101000010011010000111010110010011100101100011010100100100100000010111010101111000100100110001001001000110001110000101011100011001011000100100010000010111001001010110001110001001011000101001001101001000011101010001;
    assign base[102] = 324'b011001110011100001010100100100010010100110000010001100010110010001010111010100010100001010010111001101101000010000110110100101110001100000100101011110010101011010000010000101000011100000100001010000110101011001111001000101001001011100100011010110000110001001101000010101001001011100110001001101010111000101101000001010010100;
    assign base[103] = 324'b001001110110100101011000001100010100010110000100001100010010100101110110000100111001011001110100100000100101100100101000010001100011000101010111010000010101100010010111011000110010001101100111000100100101010010011000011001010001001001001001011110000011100010010010011100110110010101000001011101000011010110000001001001101001;
    assign base[104] = 324'b011101000110000100101001010100111000010100101001011110000011011001000001000100111000010001100101001010010111001101100100010100011000100101110010100110000101001001110110010000010011001001110001100100110100100001100101010001010011100010010001011100100110011010010010001101010111000110000100100000010111011001000010001101011001;
    assign base[105] = 324'b100100110100000100101000011001110101001001010001010001110110100000111001011001111000010110010011000100100100000110000110011101010100001110010010010000100101100000111001011101100001011110010011001001100001010001011000100001101001001100010101001001000111010100010111011001000010100110000011001101000010100110000111010100010110;
    assign base[106] = 324'b011100111001010000100001011010000101011010000100010100110111001010010001010100010010100001101001001101000111100101000101011010000011011100010010100001100011011100010010010001011001001001110001100101010100100000110110010000100110001110010101000101111000000110010111001001001000010101100011001101011000000101110110100100100100;
    assign base[107] = 324'b001001100001010010010011011110000101010101110100000100101000100101100011100100111000010101100111010000010010010001010111001000011001100000110110100000010011011001110101001010010100011010010010100000110100010101110001011101000110001110000010000101011001001100101001011101010001011001001000000110000101100101000110001100100111;
    assign base[108] = 324'b100110000110011101000101000100110010011100110101001000011001011001001000000101000010001101101000011110010101001001100011010001110001100001011001010010010001010110000010001101100111100001010111011010010011010000100001001100100100000101010111100110000110010100011000100100110110001001110100011001111001100000100100010100010011;
    assign base[109] = 324'b011110000100010100011001011000110010011010010001001001110011100001010100001101010010011010000100100101110001100100100101010000110110011100011000100000010011011110010010010001100101010001110110000101011000001010010011010101001001001100100111000110000110000101101000100101000101001100100111001000110111100001100001010101001001;
    assign base[110] = 324'b001100100101011010010111100000010100100010010100000100100101011000110111000101100111001101001000100100100101001000011000010100111001010001110110010101110110010000010010001110001001010000111001100001110110000101010010011001010010100110000001011101000011100101000001011101010011001001101000011110000011001001100100010110010001;
    assign base[111] = 324'b000100110101100001101001001001000111011001000010000101010111100110000011011110001001001001000011010100010110100100100110001110000100011101010001100001010100011100010110001110010010001101110001010110010010010001101000001010011000011001110101000100110100010100010111010000111000011000101001010001100011100100100001100001110101;
    assign base[112] = 324'b010100010110001000111000010001111001100010010111000101000110001001010011010000110010010101111001100000010110000100100011100101100101011101001000011001111000010000100001001110010101100101010100001110000111000101100010001001000001011010010011010110000111011101100101100000010010100100110100001110001001011101010100011000100001;
    assign base[113] = 324'b011100110100001001010110100000011001100000010010001110010100011101100101010101101001011100011000010000110010011001000101000100110010100101111000001100100111010010001001000101010110100110000001010101100111001001000011001001110110100001000101001110010001000101011000100101110011011000100100010010010011011000100001010110000111;
    assign base[114] = 324'b010001110110100110000011000100100101000100100101011001000111001110011000001110011000001000010101011101000110100101010011100001110001001001100100011001000001001110010010100001010111011110000010010001010110100100110001001000110111000101100100010110001001010101101001011100101000010000010011100000010100010100111001011001110010;
    assign base[115] = 324'b010000100111011000110001010110011000100100110001010001011000011001110010010110000110100100100111001101000001001001001001010101110011100000010110011000011000001001001001011100110101001101110101000110000110010000101001100001010010001100010100100101100111011101100011100010010010000101010100000110010100011101100101001010000011;
    assign base[116] = 324'b001001000011011010000001011101011001011000010101010010010111100000110010011110011000001000110101011000010100010000100111001101101001010110000001000100111001010100101000010001100111010110000110000101110100100100100011100001100001011101000011001010010101001101110010100101010110000101001000100101010100100000010010001101110110;
    assign base[117] = 324'b100110000111000101100101001100100100010001100101001000111000100100010111001100100001010010010111100001100101001000010011010101110100011010001001100010010100011000010011011101010010011101010110100110000010010000110001011001110010100001000001010110010011010101001001001100100110000101111000000100111000011101011001001001000110;
    assign base[118] = 324'b001101100101100100010111001001001000000110000010010100110100011101101001011110010100011000101000001101010001100001110001001101000110010110010010001001011001100001110001011000110100010000110110001001011001100000010111011001000111000110000101100100100011010100010011011110010010010010000110100100101000010001100011000101110101;
    assign base[119] = 324'b011010000100001101110010100101010001010110010001011001001000011100110010011100110010100100010101100001100100010001010111000110000110001100101001100001100011001001011001010000010111000100101001010000110111011010000101100101110110100000100001010101000011001100010101011101100100001010011000001001001000010110010011000101110110;
    assign base[120] = 324'b010001100101000100101001100001110011001110010111010001101000000101010010001000011000011101010011010001101001100101110011010100010100001010000110100001010110001000110111100100010100000100100100100010010110011100110101011101000010011010000101001110010001010100110001100101110010011001001000011010001001001101000001010100100111;
    assign base[121] = 324'b011000100101010010000011000101111001100010010111000100100110010000110101010000110001011110010101100001100010001010001001001100010100011101010110011101000011010101101001001000011000010100010110001001111000001110010100000101110100011001010010100110000011100101010010100000110111011001000001001101101000100101000001010100100111;
    assign base[122] = 324'b001001000001010101110110100000111001100001110110001000111001010000010101100101010011010010000001011001110010011110010101011001000011000100101000011000100100000101011000011110010011000100111000011110010010010101100100010001100111001100100101100110000001010110000010100100010111001101000110001100011001100001100100001001010111;
    assign base[123] = 324'b011000100100100100010111010110000011100101010111010010000011011000010010001110000001001001100101011101001001011101000010000101011001100000110110000101100011100000100100100101110101100010010101011100110110000100100100010000010110001110011000001001010111010101111000011001000010001110010001001000111001010101110001010001101000;
    assign base[124] = 324'b000100101001100001100111010000110101001101011000010000011001001001100111011101100100001000110101000110001001001010010101000110000100001101110110100000110001011101010110100100100100011001000111100100100011010100011000100100010110001101001000011101010010010101110011011010010010100001000001010010000010010101110001011010010011;
    assign base[125] = 324'b000101101001010010000010011100110101011100100100011000110101100010010001001110000101100100010111001001000110011001000001010100101001001101111000001010011000001101110001011001010100010100110111100001000110000100101001100001010110011110010011010000010010010001110010000101011000100101100011100100010011001001100100010110000111;
    assign base[126] = 324'b100101000111001110000010011001010001100000100101100101100001001101000111000100110110010001010111100100101000010101100010011101001000000110010011010010000001011000111001001001110101011110010011001000010101100001100100001001111000000110010100010100110110001100011001010101110110010010000010011001010100100000100011011100011001;
    assign base[127] = 324'b011101100100001000011000010100111001001100100101010010010110000101111000100010010001010101110011010001100010010000110110100110000001001001010111000101010010001101000111100010010110100101111000011001010010001100010100001001000111000100111001011010000101010110000011011101100100100100100001011000011001100000100101011101000011;

    reg [6:0] cur_seed = 7'b0;
    assign template_map = base[cur_seed];

    always @(posedge sig_new) begin
        // TODO: implement the map generator
        cur_seed <= seed[6:0];
    end
endmodule



module MaskTemplate(
    sig_new, seed,
    template_mask
);
    input sig_new;
    input [31:0] seed;
    output [80:0] template_mask;

    wire [8:0] base [31:0];
    assign base[0] = 9'b101011100;
    assign base[1] = 9'b100101100;
    assign base[2] = 9'b111100001;
    assign base[3] = 9'b100101011;
    assign base[4] = 9'b001100011;
    assign base[5] = 9'b100011010;
    assign base[6] = 9'b011100100;
    assign base[7] = 9'b101011001;
    assign base[8] = 9'b010110011;
    assign base[9] = 9'b010101010;
    assign base[10] = 9'b001011001;
    assign base[11] = 9'b001011100;
    assign base[12] = 9'b110001101;
    assign base[13] = 9'b010101110;
    assign base[14] = 9'b101101001;
    assign base[15] = 9'b010101101;
    assign base[16] = 9'b101001100;
    assign base[17] = 9'b010111010;
    assign base[18] = 9'b010001111;
    assign base[19] = 9'b111000101;
    assign base[20] = 9'b001101101;
    assign base[21] = 9'b001011011;
    assign base[22] = 9'b111000010;
    assign base[23] = 9'b011001101;
    assign base[24] = 9'b110001011;
    assign base[25] = 9'b101011001;
    assign base[26] = 9'b101100100;
    assign base[27] = 9'b101100100;
    assign base[28] = 9'b011001001;
    assign base[29] = 9'b111001001;
    assign base[30] = 9'b010011010;
    assign base[31] = 9'b111100001;

    reg [31:0] cur_seed = 32'b0;
    assign template_mask = {
        base[cur_seed[31:27]], base[cur_seed[26:22]], base[cur_seed[21:17]], base[cur_seed[16:12]],
        base[cur_seed[11:7]],
        base[cur_seed[29:25]], base[cur_seed[24:20]], base[cur_seed[19:15]], base[cur_seed[14:10]]
    };

    always @(posedge sig_new) begin
        cur_seed <= seed;
    end
endmodule